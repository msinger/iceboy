output logic [7:0] lcd_data,
output logic       n_lcd_rd,
output logic       n_lcd_wr,
output logic       n_lcd_cs,
output logic       lcd_cd,
output logic       lcd_vled,
