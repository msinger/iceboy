output logic       lcd_hsync,
output logic       lcd_vsync,
output logic       lcd_latch,
output logic       lcd_altsig,
output logic       lcd_ctrl,
output logic       lcd_clk,
output logic [1:0] lcd_data,
