.lcd_n_hsync(lcd_n_hsync_out),
.lcd_p_hsync(lcd_p_hsync_out),
.lcd_n_vsync(lcd_n_vsync_out),
.lcd_p_vsync(lcd_p_vsync_out),
.lcd_n_latch(lcd_n_latch_out),
.lcd_p_latch(lcd_p_latch_out),
.lcd_n_altsig(lcd_n_altsig_out),
.lcd_p_altsig(lcd_p_altsig_out),
.lcd_n_ctrl(lcd_n_ctrl_out),
.lcd_p_ctrl(lcd_p_ctrl_out),
.lcd_n_clk(lcd_n_clk_out),
.lcd_p_clk(lcd_p_clk_out),
.lcd_n_data(lcd_n_data_out),
.lcd_p_data(lcd_p_data_out),
